
`ifndef ETH_SEQ_PKG
`define ETH_SEQ_PKG
package eth_seq_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
import eth_env_pkg::*;
import eth_reg_pkg::*;

`include "eth_seq_lib.sv"

endpackage
`endif

