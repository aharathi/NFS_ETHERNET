`include "wishbone_package.sv"

interface wb_master_driver_if (ethmac_pif bus);

task read ();
endtask

task write();
endtask

endinterface