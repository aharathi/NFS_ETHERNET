

module hvl_top;

import uvm_pkg::*;
import eth_test_pkg::*;
initial begin 
run_test();
end 
endmodule 
